module ControleFF(
	input logic [0:8] entradas,
	output logic [0:4] saidas);